module blinky (
    input logic clk,
    input logic reset_n,
    output logic [23:0] led
);

    logic [31:0] ctr;
    assign led[23:1] = '0;

    always_ff @(posedge clk) begin
        if (~reset_n) begin
            led[0] <= '0;
            ctr <= '0;
        end
        else begin
            ctr <= ctr + 1;
            if (ctr == 12500000) begin // 12.5M = 1/2 second
                ctr <= '0;
                led[0] <= ~led[0];
            end
        end
    end

endmodule

module m_design (
    input logic clk100, // 100MHz clock
    input logic reset_n, // Active-low reset

    output logic [7:0] base_led, // LEDs on the far right side of the board
    output logic [23:0] led, // LEDs in the middle of the board

    input logic [23:0] sw, // The tiny slide-switches

    output logic [3:0] display_sel, // Select between the 4 segments
    output logic [7:0] display // Seven-segment display
);

    logic clk; // 25MHz, generated by PLL

    blinky my_blinky (
        .clk, .reset_n, .led
    );

    // 100MHz -> 25MHz
    SB_PLL40_CORE #(
//        .FEEDBACK_PATH("SIMPLE"),
//        .DIVR(4'b0000),         // DIVR =  0
//        .DIVF(7'b0000111),      // DIVF =  7
//        .DIVQ(3'b101),          // DIVQ =  5
//        .FILTER_RANGE(3'b101)   // FILTER_RANGE = 5
.FEEDBACK_PATH("SIMPLE"),
.DIVR(4'b0000),         // DIVR =  0
.DIVF(7'b0000111),      // DIVF =  7
.DIVQ(3'b100),          // DIVQ =  4
.FILTER_RANGE(3'b101)   // FILTER_RANGE = 5    
) pll (
        .LOCK(),
        .RESETB(1'b1),
        .BYPASS(1'b0),
        .REFERENCECLK(clk100),
        .PLLOUTCORE(clk)
    );

endmodule

